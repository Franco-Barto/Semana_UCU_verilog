/* Automatically generated from https://wokwi.com/projects/411379488132926465 */

`default_nettype none

// verilator lint_off UNUSEDSIGNAL
// verilator lint_off PINCONNECTEMPTY

module tt_um_wokwi_411379488132926465(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = rst_n;
  wire net2 = ui_in[0];
  wire net3 = ui_in[1];
  wire net4 = ui_in[2];
  wire net5 = ui_in[3];
  wire net6 = ui_in[4];
  wire net7 = ui_in[5];
  wire net8 = ui_in[6];
  wire net9 = ui_in[7];
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17 = 1'b1;
  wire net18 = 1'b1;
  wire net19 = 1'b0;
  wire net20 = 1'b1;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156 = 1'b0;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187 = 1'b0;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199 = 1'b1;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218 = 1'b0;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369;
  wire net370;
  wire net371;
  wire net372;
  wire net373;
  wire net374;
  wire net375;
  wire net376;
  wire net377;
  wire net378;
  wire net379;
  wire net380;
  wire net381;
  wire net382;
  wire net383;
  wire net384;
  wire net385;
  wire net386;
  wire net387;
  wire net388;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402;
  wire net403;
  wire net404;
  wire net405;
  wire net406 = 1'b0;
  wire net407;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412 = 1'b0;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421;
  wire net422;
  wire net423;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428;
  wire net429;
  wire net430;
  wire net431;
  wire net432;
  wire net433;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446;
  wire net447;
  wire net448;
  wire net449;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456;
  wire net457;
  wire net458;
  wire net459;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473;
  wire net474;
  wire net475;
  wire net476;
  wire net477;
  wire net478;
  wire net479;
  wire net480;
  wire net481;
  wire net482;
  wire net483;
  wire net484;
  wire net485;
  wire net486;
  wire net487;
  wire net488;
  wire net489;
  wire net490;
  wire net491;
  wire net492;
  wire net493;
  wire net494;
  wire net495;
  wire net496;
  wire net497;
  wire net498;
  wire net499;
  wire net500;
  wire net501;
  wire net502;
  wire net503;
  wire net504;
  wire net505;
  wire net506;
  wire net507;
  wire net508;
  wire net509;
  wire net510;
  wire net511;
  wire net512;
  wire net513;
  wire net514;
  wire net515;
  wire net516;
  wire net517;
  wire net518;
  wire net519;
  wire net520;
  wire net521 = 1'b0;
  wire net522;
  wire net523;
  wire net524;
  wire net525;
  wire net526 = 1'b1;
  wire net527 = 1'b0;
  wire net528;
  wire net529;
  wire net530;
  wire net531;
  wire net532;
  wire net533;
  wire net534;
  wire net535;
  wire net536;
  wire net537;
  wire net538;
  wire net539;
  wire net540;
  wire net541;
  wire net542;
  wire net543;
  wire net544;
  wire net545;
  wire net546;
  wire net547;
  wire net548;
  wire net549;
  wire net550;
  wire net551;
  wire net552;
  wire net553 = 1'b0;
  wire net554;
  wire net555;
  wire net556;
  wire net557;
  wire net558;
  wire net559;
  wire net560;
  wire net561;
  wire net562;
  wire net563;
  wire net564;
  wire net565;
  wire net566;
  wire net567;
  wire net568;
  wire net569;
  wire net570;
  wire net571;
  wire net572;
  wire net573;
  wire net574;
  wire net575;
  wire net576;
  wire net577;
  wire net578;
  wire net579;
  wire net580;
  wire net581;
  wire net582;
  wire net583;
  wire net584;
  wire net585;
  wire net586 = 1'b0;
  wire net587;
  wire net588;
  wire net589;
  wire net590;
  wire net591;
  wire net592;
  wire net593;
  wire net594;
  wire net595;
  wire net596;
  wire net597;
  wire net598;
  wire net599;
  wire net600;
  wire net601;
  wire net602;
  wire net603;
  wire net604;
  wire net605;
  wire net606;
  wire net607;
  wire net608;
  wire net609;
  wire net610;
  wire net611;
  wire net612;
  wire net613;
  wire net614;
  wire net615;
  wire net616;
  wire net617;

  assign uo_out[0] = net10;
  assign uo_out[1] = net11;
  assign uo_out[2] = net12;
  assign uo_out[3] = net13;
  assign uo_out[4] = net14;
  assign uo_out[5] = net15;
  assign uo_out[6] = net16;
  assign uo_out[7] = 0;
  assign uio_out[0] = 0;
  assign uio_oe[0] = 0;
  assign uio_out[1] = 0;
  assign uio_oe[1] = 0;
  assign uio_out[2] = 0;
  assign uio_oe[2] = 0;
  assign uio_out[3] = 0;
  assign uio_oe[3] = 0;
  assign uio_out[4] = 0;
  assign uio_oe[4] = 0;
  assign uio_out[5] = 0;
  assign uio_oe[5] = 0;
  assign uio_out[6] = 0;
  assign uio_oe[6] = 0;
  assign uio_out[7] = 0;
  assign uio_oe[7] = 0;

  mux_cell mux1 (
    .a (net21),
    .b (net22),
    .sel (net6),
    .out (net23)
  );
  mux_cell mux2 (
    .a (net24),
    .b (net25),
    .sel (net6),
    .out (net26)
  );
  mux_cell mux3 (
    .a (net27),
    .b (net28),
    .sel (net6),
    .out (net29)
  );
  mux_cell mux4 (
    .a (net30),
    .b (net31),
    .sel (net6),
    .out (net32)
  );
  mux_cell mux5 (
    .a (net26),
    .b (net23),
    .sel (net7),
    .out (net33)
  );
  mux_cell mux6 (
    .a (net32),
    .b (net29),
    .sel (net7),
    .out (net34)
  );
  mux_cell mux7 (
    .a (net34),
    .b (net33),
    .sel (net8),
    .out (net35)
  );
  mux_cell mux8 (
    .a (net35),
    .b (net36),
    .sel (net9),
    .out (net10)
  );
  mux_cell mux9 (
    .a (net37),
    .b (net38),
    .sel (net6),
    .out (net39)
  );
  mux_cell mux10 (
    .a (net40),
    .b (net41),
    .sel (net6),
    .out (net42)
  );
  mux_cell mux11 (
    .a (net43),
    .b (net44),
    .sel (net6),
    .out (net45)
  );
  mux_cell mux12 (
    .a (net46),
    .b (net47),
    .sel (net6),
    .out (net48)
  );
  mux_cell mux13 (
    .a (net42),
    .b (net39),
    .sel (net7),
    .out (net49)
  );
  mux_cell mux14 (
    .a (net48),
    .b (net45),
    .sel (net7),
    .out (net50)
  );
  mux_cell mux15 (
    .a (net50),
    .b (net49),
    .sel (net8),
    .out (net51)
  );
  mux_cell mux16 (
    .a (net51),
    .b (net52),
    .sel (net9),
    .out (net11)
  );
  mux_cell mux17 (
    .a (net53),
    .b (net54),
    .sel (net6),
    .out (net55)
  );
  mux_cell mux18 (
    .a (net56),
    .b (net57),
    .sel (net6),
    .out (net58)
  );
  mux_cell mux19 (
    .a (net59),
    .b (net60),
    .sel (net6),
    .out (net61)
  );
  mux_cell mux20 (
    .a (net62),
    .b (net63),
    .sel (net6),
    .out (net64)
  );
  mux_cell mux21 (
    .a (net58),
    .b (net55),
    .sel (net7),
    .out (net65)
  );
  mux_cell mux22 (
    .a (net64),
    .b (net61),
    .sel (net7),
    .out (net66)
  );
  mux_cell mux23 (
    .a (net66),
    .b (net65),
    .sel (net8),
    .out (net67)
  );
  mux_cell mux24 (
    .a (net67),
    .b (net68),
    .sel (net9),
    .out (net12)
  );
  mux_cell mux25 (
    .a (net69),
    .b (net70),
    .sel (net6),
    .out (net71)
  );
  mux_cell mux26 (
    .a (net72),
    .b (net73),
    .sel (net6),
    .out (net74)
  );
  mux_cell mux27 (
    .a (net75),
    .b (net76),
    .sel (net6),
    .out (net77)
  );
  mux_cell mux28 (
    .a (net78),
    .b (net79),
    .sel (net6),
    .out (net80)
  );
  mux_cell mux29 (
    .a (net74),
    .b (net71),
    .sel (net7),
    .out (net81)
  );
  mux_cell mux30 (
    .a (net80),
    .b (net77),
    .sel (net7),
    .out (net82)
  );
  mux_cell mux31 (
    .a (net82),
    .b (net81),
    .sel (net8),
    .out (net83)
  );
  mux_cell mux32 (
    .a (net83),
    .b (net84),
    .sel (net9),
    .out (net13)
  );
  mux_cell mux33 (
    .a (net85),
    .b (net86),
    .sel (net6),
    .out (net87)
  );
  mux_cell mux34 (
    .a (net88),
    .b (net89),
    .sel (net6),
    .out (net90)
  );
  mux_cell mux35 (
    .a (net91),
    .b (net92),
    .sel (net6),
    .out (net93)
  );
  mux_cell mux36 (
    .a (net94),
    .b (net95),
    .sel (net6),
    .out (net96)
  );
  mux_cell mux37 (
    .a (net90),
    .b (net87),
    .sel (net7),
    .out (net97)
  );
  mux_cell mux38 (
    .a (net96),
    .b (net93),
    .sel (net7),
    .out (net98)
  );
  mux_cell mux39 (
    .a (net98),
    .b (net97),
    .sel (net8),
    .out (net99)
  );
  mux_cell mux40 (
    .a (net99),
    .b (net100),
    .sel (net9),
    .out (net14)
  );
  mux_cell mux41 (
    .a (net101),
    .b (net102),
    .sel (net6),
    .out (net103)
  );
  mux_cell mux42 (
    .a (net104),
    .b (net105),
    .sel (net6),
    .out (net106)
  );
  mux_cell mux43 (
    .a (net107),
    .b (net108),
    .sel (net6),
    .out (net109)
  );
  mux_cell mux44 (
    .a (net110),
    .b (net111),
    .sel (net6),
    .out (net112)
  );
  mux_cell mux45 (
    .a (net106),
    .b (net103),
    .sel (net7),
    .out (net113)
  );
  mux_cell mux46 (
    .a (net112),
    .b (net109),
    .sel (net7),
    .out (net114)
  );
  mux_cell mux47 (
    .a (net114),
    .b (net113),
    .sel (net8),
    .out (net115)
  );
  mux_cell mux48 (
    .a (net115),
    .b (net116),
    .sel (net9),
    .out (net15)
  );
  mux_cell mux49 (
    .a (net117),
    .b (net118),
    .sel (net6),
    .out (net119)
  );
  mux_cell mux50 (
    .a (net120),
    .b (net121),
    .sel (net6),
    .out (net122)
  );
  mux_cell mux51 (
    .a (net123),
    .b (net124),
    .sel (net6),
    .out (net125)
  );
  mux_cell mux52 (
    .a (net126),
    .b (net127),
    .sel (net6),
    .out (net128)
  );
  mux_cell mux53 (
    .a (net122),
    .b (net119),
    .sel (net7),
    .out (net129)
  );
  mux_cell mux54 (
    .a (net128),
    .b (net125),
    .sel (net7),
    .out (net130)
  );
  mux_cell mux55 (
    .a (net130),
    .b (net129),
    .sel (net8),
    .out (net131)
  );
  mux_cell mux56 (
    .a (net131),
    .b (net132),
    .sel (net9),
    .out (net16)
  );
  not_cell not1 (
    .in (net3),
    .out (net133)
  );
  not_cell not2 (
    .in (net4),
    .out (net134)
  );
  not_cell not3 (
    .in (net5),
    .out (net135)
  );
  and_cell and1 (
    .a (net3),
    .b (net5),
    .out (net136)
  );
  or_cell or1 (
    .a (net136),
    .b (net137),
    .out (net138)
  );
  and_cell and2 (
    .a (net3),
    .b (net135),
    .out (net139)
  );
  and_cell and3 (
    .a (net4),
    .b (net133),
    .out (net140)
  );
  and_cell and4 (
    .a (net4),
    .b (net135),
    .out (net141)
  );
  and_cell and5 (
    .a (net3),
    .b (net134),
    .out (net142)
  );
  and_cell and6 (
    .a (net4),
    .b (net5),
    .out (net143)
  );
  and_cell and7 (
    .a (net134),
    .b (net135),
    .out (net144)
  );
  and_cell and8 (
    .a (net5),
    .b (net142),
    .out (net145)
  );
  and_cell and9 (
    .a (net133),
    .b (net135),
    .out (net137)
  );
  or_cell or2 (
    .a (net2),
    .b (net4),
    .out (net146)
  );
  or_cell or3 (
    .a (net138),
    .b (net146),
    .out (net46)
  );
  or_cell or4 (
    .a (net143),
    .b (net144),
    .out (net147)
  );
  or_cell or5 (
    .a (net147),
    .b (net133),
    .out (net30)
  );
  or_cell or6 (
    .a (net3),
    .b (net134),
    .out (net148)
  );
  or_cell or7 (
    .a (net148),
    .b (net5),
    .out (net126)
  );
  or_cell or8 (
    .a (net141),
    .b (net140),
    .out (net149)
  );
  or_cell or9 (
    .a (net2),
    .b (net137),
    .out (net150)
  );
  or_cell or10 (
    .a (net149),
    .b (net150),
    .out (net151)
  );
  or_cell or11 (
    .a (net151),
    .b (net145),
    .out (net110)
  );
  or_cell or12 (
    .a (net141),
    .b (net137),
    .out (net94)
  );
  or_cell or13 (
    .a (net142),
    .b (net139),
    .out (net152)
  );
  or_cell or14 (
    .a (net144),
    .b (net2),
    .out (net153)
  );
  or_cell or15 (
    .a (net152),
    .b (net153),
    .out (net62)
  );
  or_cell or16 (
    .a (net141),
    .b (net142),
    .out (net154)
  );
  or_cell or17 (
    .a (net2),
    .b (net140),
    .out (net155)
  );
  or_cell or18 (
    .a (net154),
    .b (net155),
    .out (net78)
  );
  not_cell not4 (
    .in (net157),
    .out (net158)
  );
  not_cell not5 (
    .in (net159),
    .out (net160)
  );
  not_cell not6 (
    .in (net161),
    .out (net162)
  );
  and_cell and10 (
    .a (net159),
    .b (net157),
    .out (net163)
  );
  and_cell and11 (
    .a (net161),
    .b (net158),
    .out (net164)
  );
  and_cell and12 (
    .a (net159),
    .b (net158),
    .out (net165)
  );
  and_cell and13 (
    .a (net160),
    .b (net158),
    .out (net166)
  );
  and_cell and14 (
    .a (net162),
    .b (net158),
    .out (net167)
  );
  and_cell and15 (
    .a (net161),
    .b (net157),
    .out (net168)
  );
  and_cell and16 (
    .a (net159),
    .b (net162),
    .out (net169)
  );
  and_cell and17 (
    .a (net160),
    .b (net161),
    .out (net170)
  );
  and_cell and18 (
    .a (net159),
    .b (net162),
    .out (net171)
  );
  or_cell or19 (
    .a (net172),
    .b (net173),
    .out (net31)
  );
  or_cell or20 (
    .a (net163),
    .b (net161),
    .out (net173)
  );
  or_cell or21 (
    .a (net174),
    .b (net166),
    .out (net172)
  );
  or_cell or22 (
    .a (net175),
    .b (net176),
    .out (net47)
  );
  or_cell or23 (
    .a (net168),
    .b (net167),
    .out (net176)
  );
  or_cell or24 (
    .a (net160),
    .b (net174),
    .out (net175)
  );
  or_cell or25 (
    .a (net164),
    .b (net170),
    .out (net177)
  );
  or_cell or26 (
    .a (net178),
    .b (net157),
    .out (net63)
  );
  or_cell or27 (
    .a (net159),
    .b (net167),
    .out (net178)
  );
  or_cell or28 (
    .a (net177),
    .b (net179),
    .out (net79)
  );
  or_cell or29 (
    .a (net166),
    .b (net180),
    .out (net179)
  );
  and_cell and19 (
    .a (net158),
    .b (net181),
    .out (net95)
  );
  not_cell not7 (
    .in (net169),
    .out (net181)
  );
  or_cell or30 (
    .a (net182),
    .b (net183),
    .out (net111)
  );
  or_cell or31 (
    .a (net167),
    .b (net169),
    .out (net183)
  );
  or_cell or32 (
    .a (net174),
    .b (net165),
    .out (net182)
  );
  or_cell or33 (
    .a (net184),
    .b (net185),
    .out (net127)
  );
  or_cell or34 (
    .a (net170),
    .b (net169),
    .out (net185)
  );
  or_cell or35 (
    .a (net174),
    .b (net164),
    .out (net184)
  );
  and_cell and20 (
    .a (net171),
    .b (net157),
    .out (net180)
  );
  dffsr_cell flop1 (
    .d (net186),
    .clk (net2),
    .s (net187),
    .r (net188),
    .q (net157),
    .notq (net189)
  );
  dffsr_cell flop2 (
    .d (net190),
    .clk (net2),
    .s (net187),
    .r (net188),
    .q (net161),
    .notq (net191)
  );
  dffsr_cell flop3 (
    .d (net192),
    .clk (net2),
    .s (net187),
    .r (net188),
    .q (net174),
    .notq (net193)
  );
  dffsr_cell flop4 (
    .d (net194),
    .clk (net2),
    .s (net187),
    .r (net188),
    .q (net159),
    .notq (net195)
  );
  not_cell not8 (
    .in (net1),
    .out (net188)
  );
  and_cell and21 (
    .a (net191),
    .b (net157),
    .out (net196)
  );
  and_cell and22 (
    .a (net174),
    .b (net195),
    .out (net197)
  );
  and_cell and23 (
    .a (net196),
    .b (net197),
    .out (net198)
  );
  or_cell or36 (
    .a (net200),
    .b (net201),
    .out (net202)
  );
  and_cell and24 (
    .a (net189),
    .b (net199),
    .out (net200)
  );
  and_cell and25 (
    .a (net203),
    .b (net157),
    .out (net201)
  );
  not_cell not9 (
    .in (net199),
    .out (net203)
  );
  and_cell and26 (
    .a (net204),
    .b (net202),
    .out (net186)
  );
  not_cell not10 (
    .in (net198),
    .out (net204)
  );
  and_cell and27 (
    .a (net191),
    .b (net157),
    .out (net205)
  );
  and_cell and28 (
    .a (net206),
    .b (net161),
    .out (net207)
  );
  not_cell not11 (
    .in (net157),
    .out (net206)
  );
  or_cell or37 (
    .a (net205),
    .b (net207),
    .out (net208)
  );
  or_cell or38 (
    .a (net209),
    .b (net210),
    .out (net194)
  );
  and_cell and29 (
    .a (net195),
    .b (net211),
    .out (net209)
  );
  and_cell and30 (
    .a (net212),
    .b (net159),
    .out (net210)
  );
  not_cell not12 (
    .in (net211),
    .out (net212)
  );
  and_cell and31 (
    .a (net157),
    .b (net161),
    .out (net211)
  );
  or_cell or39 (
    .a (net213),
    .b (net214),
    .out (net215)
  );
  and_cell and32 (
    .a (net193),
    .b (net216),
    .out (net213)
  );
  and_cell and33 (
    .a (net217),
    .b (net174),
    .out (net214)
  );
  not_cell not13 (
    .in (net216),
    .out (net217)
  );
  and_cell and34 (
    .a (net159),
    .b (net211),
    .out (net216)
  );
  and_cell and35 (
    .a (net215),
    .b (net204),
    .out (net192)
  );
  and_cell and36 (
    .a (net208),
    .b (net204),
    .out (net190)
  );
  and_cell and37 (
    .a (net219),
    .b (net220),
    .out (net221)
  );
  and_cell and38 (
    .a (net2),
    .b (net4),
    .out (net222)
  );
  or_cell or40 (
    .a (net221),
    .b (net222),
    .out (net223)
  );
  or_cell or41 (
    .a (net223),
    .b (net3),
    .out (net27)
  );
  not_cell not14 (
    .in (net2),
    .out (net219)
  );
  not_cell not15 (
    .in (net4),
    .out (net220)
  );
  and_cell and39 (
    .a (net224),
    .b (net225),
    .out (net226)
  );
  and_cell and40 (
    .a (net3),
    .b (net4),
    .out (net227)
  );
  or_cell or42 (
    .a (net226),
    .b (net227),
    .out (net228)
  );
  or_cell or43 (
    .a (net228),
    .b (net229),
    .out (net43)
  );
  not_cell not16 (
    .in (net3),
    .out (net224)
  );
  not_cell not17 (
    .in (net4),
    .out (net225)
  );
  not_cell not18 (
    .in (net2),
    .out (net229)
  );
  or_cell or44 (
    .a (net230),
    .b (net4),
    .out (net231)
  );
  or_cell or45 (
    .a (net231),
    .b (net2),
    .out (net59)
  );
  not_cell not19 (
    .in (net3),
    .out (net230)
  );
  and_cell and41 (
    .a (net232),
    .b (net233),
    .out (net234)
  );
  and_cell and42 (
    .a (net232),
    .b (net3),
    .out (net235)
  );
  and_cell and43 (
    .a (net236),
    .b (net4),
    .out (net237)
  );
  and_cell and44 (
    .a (net3),
    .b (net238),
    .out (net239)
  );
  or_cell or46 (
    .a (net234),
    .b (net235),
    .out (net240)
  );
  or_cell or47 (
    .a (net240),
    .b (net241),
    .out (net75)
  );
  or_cell or48 (
    .a (net237),
    .b (net239),
    .out (net241)
  );
  and_cell and45 (
    .a (net2),
    .b (net242),
    .out (net236)
  );
  not_cell not20 (
    .in (net2),
    .out (net232)
  );
  not_cell not21 (
    .in (net4),
    .out (net233)
  );
  not_cell not22 (
    .in (net3),
    .out (net242)
  );
  not_cell not23 (
    .in (net4),
    .out (net238)
  );
  and_cell and46 (
    .a (net243),
    .b (net244),
    .out (net245)
  );
  and_cell and47 (
    .a (net3),
    .b (net246),
    .out (net247)
  );
  or_cell or49 (
    .a (net245),
    .b (net247),
    .out (net91)
  );
  not_cell not24 (
    .in (net2),
    .out (net243)
  );
  not_cell not25 (
    .in (net4),
    .out (net244)
  );
  not_cell not26 (
    .in (net4),
    .out (net246)
  );
  and_cell and48 (
    .a (net248),
    .b (net249),
    .out (net250)
  );
  and_cell and49 (
    .a (net2),
    .b (net251),
    .out (net252)
  );
  and_cell and50 (
    .a (net2),
    .b (net253),
    .out (net254)
  );
  or_cell or50 (
    .a (net250),
    .b (net252),
    .out (net255)
  );
  or_cell or51 (
    .a (net255),
    .b (net254),
    .out (net107)
  );
  not_cell not27 (
    .in (net3),
    .out (net248)
  );
  not_cell not28 (
    .in (net4),
    .out (net249)
  );
  not_cell not29 (
    .in (net3),
    .out (net251)
  );
  not_cell not30 (
    .in (net4),
    .out (net253)
  );
  and_cell and51 (
    .a (net256),
    .b (net3),
    .out (net257)
  );
  and_cell and52 (
    .a (net2),
    .b (net258),
    .out (net259)
  );
  and_cell and53 (
    .a (net3),
    .b (net260),
    .out (net261)
  );
  or_cell or52 (
    .a (net257),
    .b (net259),
    .out (net262)
  );
  or_cell or53 (
    .a (net262),
    .b (net261),
    .out (net123)
  );
  not_cell not31 (
    .in (net2),
    .out (net256)
  );
  not_cell not32 (
    .in (net3),
    .out (net258)
  );
  not_cell not33 (
    .in (net4),
    .out (net260)
  );
  and_cell and54 (
    .a (net263),
    .b (net264),
    .out (net265)
  );
  not_cell not34 (
    .in (net2),
    .out (net263)
  );
  or_cell or54 (
    .a (net3),
    .b (net265),
    .out (net266)
  );
  or_cell or55 (
    .a (net266),
    .b (net267),
    .out (net28)
  );
  and_cell and55 (
    .a (net2),
    .b (net4),
    .out (net267)
  );
  not_cell not35 (
    .in (net4),
    .out (net264)
  );
  or_cell or56 (
    .a (net268),
    .b (net269),
    .out (net44)
  );
  or_cell or57 (
    .a (net270),
    .b (net271),
    .out (net268)
  );
  and_cell and56 (
    .a (net3),
    .b (net4),
    .out (net269)
  );
  and_cell and57 (
    .a (net272),
    .b (net273),
    .out (net271)
  );
  not_cell not36 (
    .in (net4),
    .out (net273)
  );
  not_cell not37 (
    .in (net3),
    .out (net272)
  );
  not_cell not38 (
    .in (net2),
    .out (net270)
  );
  or_cell or58 (
    .a (net274),
    .b (net275),
    .out (net60)
  );
  or_cell or59 (
    .a (net2),
    .b (net4),
    .out (net274)
  );
  not_cell not39 (
    .in (net3),
    .out (net275)
  );
  or_cell or60 (
    .a (net276),
    .b (net277),
    .out (net278)
  );
  or_cell or61 (
    .a (net279),
    .b (net280),
    .out (net281)
  );
  or_cell or62 (
    .a (net278),
    .b (net281),
    .out (net76)
  );
  and_cell and58 (
    .a (net282),
    .b (net283),
    .out (net276)
  );
  and_cell and59 (
    .a (net284),
    .b (net3),
    .out (net277)
  );
  not_cell not40 (
    .in (net2),
    .out (net284)
  );
  not_cell not41 (
    .in (net4),
    .out (net283)
  );
  not_cell not42 (
    .in (net2),
    .out (net282)
  );
  not_cell not43 (
    .in (net3),
    .out (net285)
  );
  not_cell not44 (
    .in (net2),
    .out (net286)
  );
  and_cell and60 (
    .a (net2),
    .b (net287),
    .out (net280)
  );
  and_cell and61 (
    .a (net3),
    .b (net288),
    .out (net279)
  );
  and_cell and62 (
    .a (net285),
    .b (net4),
    .out (net287)
  );
  or_cell or63 (
    .a (net289),
    .b (net290),
    .out (net92)
  );
  and_cell and63 (
    .a (net286),
    .b (net291),
    .out (net289)
  );
  and_cell and64 (
    .a (net3),
    .b (net292),
    .out (net290)
  );
  not_cell not45 (
    .in (net4),
    .out (net292)
  );
  not_cell not46 (
    .in (net4),
    .out (net291)
  );
  or_cell or64 (
    .a (net293),
    .b (net294),
    .out (net108)
  );
  or_cell or65 (
    .a (net295),
    .b (net296),
    .out (net293)
  );
  and_cell and65 (
    .a (net297),
    .b (net298),
    .out (net295)
  );
  and_cell and66 (
    .a (net2),
    .b (net299),
    .out (net296)
  );
  and_cell and67 (
    .a (net2),
    .b (net300),
    .out (net294)
  );
  not_cell not47 (
    .in (net4),
    .out (net300)
  );
  not_cell not48 (
    .in (net3),
    .out (net297)
  );
  not_cell not49 (
    .in (net3),
    .out (net299)
  );
  not_cell not50 (
    .in (net4),
    .out (net298)
  );
  or_cell or66 (
    .a (net301),
    .b (net302),
    .out (net124)
  );
  or_cell or67 (
    .a (net303),
    .b (net304),
    .out (net301)
  );
  and_cell and68 (
    .a (net2),
    .b (net305),
    .out (net302)
  );
  and_cell and69 (
    .a (net3),
    .b (net306),
    .out (net304)
  );
  and_cell and70 (
    .a (net307),
    .b (net3),
    .out (net303)
  );
  not_cell not51 (
    .in (net2),
    .out (net307)
  );
  not_cell not52 (
    .in (net3),
    .out (net305)
  );
  not_cell not53 (
    .in (net4),
    .out (net306)
  );
  not_cell not54 (
    .in (net4),
    .out (net288)
  );
  and_cell and71 (
    .a (net2),
    .b (net308),
    .out (net309)
  );
  not_cell not55 (
    .in (net3),
    .out (net308)
  );
  or_cell or68 (
    .a (net310),
    .b (net311),
    .out (net104)
  );
  or_cell or69 (
    .a (net309),
    .b (net312),
    .out (net310)
  );
  and_cell and72 (
    .a (net2),
    .b (net313),
    .out (net312)
  );
  and_cell and73 (
    .a (net314),
    .b (net315),
    .out (net311)
  );
  not_cell not56 (
    .in (net4),
    .out (net313)
  );
  not_cell not57 (
    .in (net4),
    .out (net315)
  );
  not_cell not58 (
    .in (net3),
    .out (net314)
  );
  and_cell and74 (
    .a (net316),
    .b (net2),
    .out (net317)
  );
  not_cell not59 (
    .in (net3),
    .out (net316)
  );
  or_cell or70 (
    .a (net317),
    .b (net318),
    .out (net319)
  );
  and_cell and75 (
    .a (net2),
    .b (net320),
    .out (net318)
  );
  not_cell not60 (
    .in (net4),
    .out (net320)
  );
  or_cell or71 (
    .a (net319),
    .b (net321),
    .out (net120)
  );
  and_cell and76 (
    .a (net322),
    .b (net3),
    .out (net321)
  );
  not_cell not61 (
    .in (net2),
    .out (net322)
  );
  not_cell not62 (
    .in (net4),
    .out (net323)
  );
  and_cell and77 (
    .a (net323),
    .b (net3),
    .out (net324)
  );
  or_cell or72 (
    .a (net324),
    .b (net325),
    .out (net88)
  );
  not_cell not63 (
    .in (net4),
    .out (net326)
  );
  not_cell not64 (
    .in (net2),
    .out (net327)
  );
  and_cell and78 (
    .a (net327),
    .b (net326),
    .out (net325)
  );
  or_cell or73 (
    .a (net2),
    .b (net4),
    .out (net328)
  );
  or_cell or74 (
    .a (net328),
    .b (net329),
    .out (net56)
  );
  not_cell not65 (
    .in (net3),
    .out (net329)
  );
  not_cell not66 (
    .in (net4),
    .out (net330)
  );
  not_cell not67 (
    .in (net2),
    .out (net331)
  );
  or_cell or75 (
    .a (net332),
    .b (net333),
    .out (net334)
  );
  and_cell and79 (
    .a (net331),
    .b (net330),
    .out (net332)
  );
  and_cell and80 (
    .a (net335),
    .b (net3),
    .out (net333)
  );
  not_cell not68 (
    .in (net2),
    .out (net335)
  );
  not_cell not69 (
    .in (net4),
    .out (net336)
  );
  and_cell and81 (
    .a (net336),
    .b (net3),
    .out (net337)
  );
  and_cell and82 (
    .a (net2),
    .b (net4),
    .out (net338)
  );
  and_cell and83 (
    .a (net338),
    .b (net339),
    .out (net340)
  );
  not_cell not70 (
    .in (net3),
    .out (net339)
  );
  or_cell or76 (
    .a (net337),
    .b (net340),
    .out (net341)
  );
  or_cell or77 (
    .a (net334),
    .b (net341),
    .out (net72)
  );
  or_cell or78 (
    .a (net342),
    .b (net343),
    .out (net344)
  );
  not_cell not71 (
    .in (net2),
    .out (net345)
  );
  not_cell not72 (
    .in (net2),
    .out (net346)
  );
  and_cell and84 (
    .a (net345),
    .b (net347),
    .out (net342)
  );
  and_cell and85 (
    .a (net346),
    .b (net3),
    .out (net343)
  );
  or_cell or79 (
    .a (net344),
    .b (net348),
    .out (net24)
  );
  and_cell and86 (
    .a (net2),
    .b (net4),
    .out (net348)
  );
  not_cell not73 (
    .in (net4),
    .out (net347)
  );
  not_cell not74 (
    .in (net2),
    .out (net349)
  );
  not_cell not75 (
    .in (net3),
    .out (net350)
  );
  not_cell not76 (
    .in (net4),
    .out (net351)
  );
  and_cell and87 (
    .a (net350),
    .b (net351),
    .out (net352)
  );
  or_cell or80 (
    .a (net353),
    .b (net354),
    .out (net40)
  );
  or_cell or81 (
    .a (net349),
    .b (net352),
    .out (net353)
  );
  and_cell and88 (
    .a (net3),
    .b (net4),
    .out (net354)
  );
  or_cell or82 (
    .a (net355),
    .b (net356),
    .out (net357)
  );
  not_cell not77 (
    .in (net358),
    .out (net359)
  );
  not_cell not78 (
    .in (net360),
    .out (net361)
  );
  not_cell not79 (
    .in (net360),
    .out (net362)
  );
  and_cell and89 (
    .a (net361),
    .b (net359),
    .out (net355)
  );
  and_cell and90 (
    .a (net362),
    .b (net363),
    .out (net356)
  );
  or_cell or83 (
    .a (net357),
    .b (net364),
    .out (net25)
  );
  and_cell and91 (
    .a (net360),
    .b (net358),
    .out (net364)
  );
  not_cell not80 (
    .in (net360),
    .out (net365)
  );
  not_cell not81 (
    .in (net363),
    .out (net366)
  );
  not_cell not82 (
    .in (net358),
    .out (net367)
  );
  and_cell and92 (
    .a (net366),
    .b (net367),
    .out (net368)
  );
  or_cell or84 (
    .a (net369),
    .b (net370),
    .out (net41)
  );
  or_cell or85 (
    .a (net365),
    .b (net368),
    .out (net369)
  );
  and_cell and93 (
    .a (net363),
    .b (net358),
    .out (net370)
  );
  or_cell or86 (
    .a (net360),
    .b (net358),
    .out (net371)
  );
  or_cell or87 (
    .a (net371),
    .b (net372),
    .out (net57)
  );
  not_cell not83 (
    .in (net363),
    .out (net372)
  );
  not_cell not84 (
    .in (net358),
    .out (net373)
  );
  not_cell not85 (
    .in (net360),
    .out (net374)
  );
  or_cell or88 (
    .a (net375),
    .b (net376),
    .out (net377)
  );
  and_cell and94 (
    .a (net374),
    .b (net373),
    .out (net375)
  );
  and_cell and95 (
    .a (net378),
    .b (net363),
    .out (net376)
  );
  not_cell not86 (
    .in (net360),
    .out (net378)
  );
  not_cell not87 (
    .in (net358),
    .out (net379)
  );
  and_cell and96 (
    .a (net379),
    .b (net363),
    .out (net380)
  );
  and_cell and97 (
    .a (net360),
    .b (net358),
    .out (net381)
  );
  and_cell and98 (
    .a (net381),
    .b (net382),
    .out (net383)
  );
  not_cell not88 (
    .in (net363),
    .out (net382)
  );
  or_cell or89 (
    .a (net380),
    .b (net383),
    .out (net384)
  );
  or_cell or90 (
    .a (net377),
    .b (net384),
    .out (net73)
  );
  not_cell not89 (
    .in (net358),
    .out (net385)
  );
  and_cell and99 (
    .a (net385),
    .b (net363),
    .out (net386)
  );
  or_cell or91 (
    .a (net386),
    .b (net387),
    .out (net89)
  );
  not_cell not90 (
    .in (net358),
    .out (net388)
  );
  not_cell not91 (
    .in (net360),
    .out (net389)
  );
  and_cell and100 (
    .a (net389),
    .b (net388),
    .out (net387)
  );
  and_cell and101 (
    .a (net360),
    .b (net390),
    .out (net391)
  );
  not_cell not92 (
    .in (net363),
    .out (net390)
  );
  or_cell or92 (
    .a (net392),
    .b (net393),
    .out (net105)
  );
  or_cell or93 (
    .a (net391),
    .b (net394),
    .out (net392)
  );
  and_cell and102 (
    .a (net360),
    .b (net395),
    .out (net394)
  );
  and_cell and103 (
    .a (net396),
    .b (net397),
    .out (net393)
  );
  not_cell not93 (
    .in (net358),
    .out (net395)
  );
  not_cell not94 (
    .in (net358),
    .out (net397)
  );
  not_cell not95 (
    .in (net363),
    .out (net396)
  );
  and_cell and104 (
    .a (net398),
    .b (net360),
    .out (net399)
  );
  not_cell not96 (
    .in (net363),
    .out (net398)
  );
  or_cell or94 (
    .a (net399),
    .b (net400),
    .out (net401)
  );
  and_cell and105 (
    .a (net360),
    .b (net402),
    .out (net400)
  );
  not_cell not97 (
    .in (net358),
    .out (net402)
  );
  or_cell or95 (
    .a (net401),
    .b (net403),
    .out (net121)
  );
  and_cell and106 (
    .a (net404),
    .b (net363),
    .out (net403)
  );
  not_cell not98 (
    .in (net360),
    .out (net404)
  );
  dffsr_cell flop5 (
    .d (net405),
    .clk (net2),
    .s (net406),
    .r (net407),
    .q (net358),
    .notq (net405)
  );
  dffsr_cell flop6 (
    .d (net408),
    .clk (net405),
    .s (net406),
    .r (net407),
    .q (net363),
    .notq (net408)
  );
  dffsr_cell flop7 (
    .d (net409),
    .clk (net408),
    .s (net406),
    .r (net407),
    .q (net360),
    .notq (net409)
  );
  not_cell not99 (
    .in (net1),
    .out (net407)
  );
  dffsr_cell flop8 (
    .d (net410),
    .clk (net411),
    .s (net412),
    .r (net413),
    .q (net414),
    .notq (net410)
  );
  dffsr_cell flop9 (
    .d (net411),
    .clk (net415),
    .s (net412),
    .r (net413),
    .q (net416),
    .notq (net411)
  );
  dffsr_cell flop10 (
    .d (net415),
    .clk (net417),
    .s (net412),
    .r (net413),
    .q (net418),
    .notq (net415)
  );
  dffsr_cell flop11 (
    .d (net417),
    .clk (net2),
    .s (net412),
    .r (net413),
    .q (net419),
    .notq (net417)
  );
  not_cell not100 (
    .in (net1),
    .out (net413)
  );
  not_cell not101 (
    .in (net416),
    .out (net420)
  );
  not_cell not102 (
    .in (net418),
    .out (net421)
  );
  not_cell not103 (
    .in (net419),
    .out (net422)
  );
  and_cell and107 (
    .a (net416),
    .b (net419),
    .out (net423)
  );
  or_cell or96 (
    .a (net423),
    .b (net424),
    .out (net425)
  );
  and_cell and108 (
    .a (net416),
    .b (net422),
    .out (net426)
  );
  and_cell and109 (
    .a (net418),
    .b (net420),
    .out (net427)
  );
  and_cell and110 (
    .a (net418),
    .b (net422),
    .out (net428)
  );
  and_cell and111 (
    .a (net416),
    .b (net421),
    .out (net429)
  );
  and_cell and112 (
    .a (net418),
    .b (net419),
    .out (net430)
  );
  and_cell and113 (
    .a (net421),
    .b (net422),
    .out (net431)
  );
  and_cell and114 (
    .a (net419),
    .b (net429),
    .out (net432)
  );
  and_cell and115 (
    .a (net420),
    .b (net422),
    .out (net424)
  );
  or_cell or97 (
    .a (net414),
    .b (net418),
    .out (net433)
  );
  or_cell or98 (
    .a (net425),
    .b (net433),
    .out (net21)
  );
  or_cell or99 (
    .a (net430),
    .b (net431),
    .out (net434)
  );
  or_cell or100 (
    .a (net434),
    .b (net420),
    .out (net37)
  );
  or_cell or101 (
    .a (net416),
    .b (net421),
    .out (net435)
  );
  or_cell or102 (
    .a (net435),
    .b (net419),
    .out (net53)
  );
  or_cell or103 (
    .a (net428),
    .b (net427),
    .out (net436)
  );
  or_cell or104 (
    .a (net414),
    .b (net424),
    .out (net437)
  );
  or_cell or105 (
    .a (net436),
    .b (net437),
    .out (net438)
  );
  or_cell or106 (
    .a (net438),
    .b (net432),
    .out (net69)
  );
  or_cell or107 (
    .a (net428),
    .b (net424),
    .out (net85)
  );
  or_cell or108 (
    .a (net429),
    .b (net426),
    .out (net439)
  );
  or_cell or109 (
    .a (net431),
    .b (net414),
    .out (net440)
  );
  or_cell or110 (
    .a (net439),
    .b (net440),
    .out (net101)
  );
  or_cell or111 (
    .a (net428),
    .b (net429),
    .out (net441)
  );
  or_cell or112 (
    .a (net414),
    .b (net427),
    .out (net442)
  );
  or_cell or113 (
    .a (net441),
    .b (net442),
    .out (net117)
  );
  not_cell not104 (
    .in (net1),
    .out (net443)
  );
  not_cell not105 (
    .in (net444),
    .out (net445)
  );
  not_cell not106 (
    .in (net446),
    .out (net447)
  );
  not_cell not107 (
    .in (net448),
    .out (net449)
  );
  and_cell and116 (
    .a (net448),
    .b (net446),
    .out (net450)
  );
  and_cell and117 (
    .a (net449),
    .b (net447),
    .out (net451)
  );
  or_cell or114 (
    .a (net450),
    .b (net444),
    .out (net452)
  );
  or_cell or115 (
    .a (net452),
    .b (net451),
    .out (net453)
  );
  or_cell or116 (
    .a (net447),
    .b (net454),
    .out (net455)
  );
  and_cell and118 (
    .a (net448),
    .b (net444),
    .out (net454)
  );
  and_cell and119 (
    .a (net449),
    .b (net445),
    .out (net456)
  );
  or_cell or117 (
    .a (net455),
    .b (net456),
    .out (net457)
  );
  or_cell or118 (
    .a (net448),
    .b (net446),
    .out (net458)
  );
  or_cell or119 (
    .a (net458),
    .b (net445),
    .out (net459)
  );
  or_cell or120 (
    .a (net460),
    .b (net461),
    .out (net462)
  );
  and_cell and120 (
    .a (net444),
    .b (net447),
    .out (net460)
  );
  and_cell and121 (
    .a (net449),
    .b (net444),
    .out (net461)
  );
  and_cell and122 (
    .a (net449),
    .b (net447),
    .out (net463)
  );
  and_cell and123 (
    .a (net448),
    .b (net446),
    .out (net464)
  );
  and_cell and124 (
    .a (net464),
    .b (net445),
    .out (net465)
  );
  or_cell or121 (
    .a (net463),
    .b (net465),
    .out (net466)
  );
  or_cell or122 (
    .a (net462),
    .b (net466),
    .out (net467)
  );
  or_cell or123 (
    .a (net468),
    .b (net469),
    .out (net470)
  );
  and_cell and125 (
    .a (net449),
    .b (net444),
    .out (net468)
  );
  and_cell and126 (
    .a (net449),
    .b (net447),
    .out (net469)
  );
  and_cell and127 (
    .a (net446),
    .b (net445),
    .out (net471)
  );
  or_cell or124 (
    .a (net471),
    .b (net472),
    .out (net473)
  );
  and_cell and128 (
    .a (net449),
    .b (net446),
    .out (net472)
  );
  and_cell and129 (
    .a (net449),
    .b (net445),
    .out (net474)
  );
  or_cell or125 (
    .a (net473),
    .b (net474),
    .out (net475)
  );
  and_cell and130 (
    .a (net446),
    .b (net445),
    .out (net476)
  );
  and_cell and131 (
    .a (net449),
    .b (net446),
    .out (net477)
  );
  or_cell or126 (
    .a (net476),
    .b (net477),
    .out (net478)
  );
  and_cell and132 (
    .a (net447),
    .b (net444),
    .out (net479)
  );
  or_cell or127 (
    .a (net478),
    .b (net479),
    .out (net480)
  );
  not_cell not108 (
    .in (net453),
    .out (net22)
  );
  not_cell not109 (
    .in (net457),
    .out (net38)
  );
  not_cell not110 (
    .in (net467),
    .out (net70)
  );
  not_cell not111 (
    .in (net459),
    .out (net54)
  );
  not_cell not112 (
    .in (net480),
    .out (net118)
  );
  not_cell not113 (
    .in (net475),
    .out (net102)
  );
  not_cell not114 (
    .in (net470),
    .out (net86)
  );
  dffsr_cell flop12 (
    .d (net481),
    .clk (net3),
    .s (net2),
    .r (net443),
    .q (net448),
    .notq (net481)
  );
  dffsr_cell flop13 (
    .d (net482),
    .clk (net483),
    .s (net2),
    .r (net443),
    .q (net446),
    .notq (net482)
  );
  dffsr_cell flop14 (
    .d (net483),
    .clk (net481),
    .s (net2),
    .r (net443),
    .q (net444),
    .notq (net483)
  );
  not_cell not115 (
    .in (net484),
    .out (net485)
  );
  not_cell not116 (
    .in (net486),
    .out (net487)
  );
  not_cell not117 (
    .in (net488),
    .out (net489)
  );
  and_cell and133 (
    .a (net487),
    .b (net489),
    .out (net490)
  );
  and_cell and134 (
    .a (net486),
    .b (net488),
    .out (net491)
  );
  and_cell and135 (
    .a (net487),
    .b (net484),
    .out (net492)
  );
  and_cell and136 (
    .a (net493),
    .b (net485),
    .out (net494)
  );
  and_cell and137 (
    .a (net486),
    .b (net488),
    .out (net493)
  );
  and_cell and138 (
    .a (net484),
    .b (net489),
    .out (net495)
  );
  and_cell and139 (
    .a (net485),
    .b (net489),
    .out (net496)
  );
  and_cell and140 (
    .a (net484),
    .b (net488),
    .out (net497)
  );
  and_cell and141 (
    .a (net486),
    .b (net489),
    .out (net498)
  );
  and_cell and142 (
    .a (net486),
    .b (net485),
    .out (net499)
  );
  or_cell or128 (
    .a (net500),
    .b (net501),
    .out (net502)
  );
  or_cell or129 (
    .a (net503),
    .b (net504),
    .out (net505)
  );
  or_cell or130 (
    .a (net506),
    .b (net507),
    .out (net508)
  );
  or_cell or131 (
    .a (net490),
    .b (net495),
    .out (net509)
  );
  or_cell or132 (
    .a (net510),
    .b (net496),
    .out (net511)
  );
  or_cell or133 (
    .a (net512),
    .b (net513),
    .out (net514)
  );
  or_cell or134 (
    .a (net496),
    .b (net499),
    .out (net503)
  );
  or_cell or135 (
    .a (net515),
    .b (net498),
    .out (net504)
  );
  or_cell or136 (
    .a (net516),
    .b (net492),
    .out (net517)
  );
  or_cell or137 (
    .a (net518),
    .b (net519),
    .out (net516)
  );
  or_cell or138 (
    .a (net495),
    .b (net494),
    .out (net519)
  );
  or_cell or139 (
    .a (net515),
    .b (net490),
    .out (net518)
  );
  or_cell or140 (
    .a (net486),
    .b (net488),
    .out (net510)
  );
  or_cell or141 (
    .a (net497),
    .b (net496),
    .out (net513)
  );
  or_cell or142 (
    .a (net515),
    .b (net487),
    .out (net512)
  );
  or_cell or143 (
    .a (net491),
    .b (net484),
    .out (net501)
  );
  or_cell or144 (
    .a (net515),
    .b (net490),
    .out (net500)
  );
  or_cell or145 (
    .a (net515),
    .b (net499),
    .out (net506)
  );
  or_cell or146 (
    .a (net498),
    .b (net492),
    .out (net507)
  );
  not_cell not118 (
    .in (net1),
    .out (net520)
  );
  dffsr_cell flop15 (
    .d (net522),
    .clk (net523),
    .s (net521),
    .r (net520),
    .q (net484),
    .notq (net522)
  );
  dffsr_cell flop16 (
    .d (net524),
    .clk (net522),
    .s (net521),
    .r (net520),
    .q (net486),
    .notq (net524)
  );
  dffsr_cell flop17 (
    .d (net523),
    .clk (net2),
    .s (net521),
    .r (net520),
    .q (net488),
    .notq (net523)
  );
  dffsr_cell flop18 (
    .d (net525),
    .clk (net524),
    .s (net521),
    .r (net520),
    .q (net515),
    .notq (net525)
  );
  dffsr_cell flop19 (
    .d (net2),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net529),
    .notq (net530)
  );
  dffsr_cell flop20 (
    .d (net529),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net531),
    .notq (net532)
  );
  dffsr_cell flop21 (
    .d (net531),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net533),
    .notq (net534)
  );
  dffsr_cell flop22 (
    .d (net533),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net535),
    .notq (net536)
  );
  dffsr_cell flop23 (
    .d (net535),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net537),
    .notq (net538)
  );
  dffsr_cell flop24 (
    .d (net537),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net539),
    .notq (net540)
  );
  dffsr_cell flop25 (
    .d (net539),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net541),
    .notq (net542)
  );
  dffsr_cell flop26 (
    .d (net541),
    .clk (net3),
    .s (net527),
    .r (net528),
    .q (net543),
    .notq ()
  );
  not_cell not119 (
    .in (net1),
    .out (net528)
  );
  mux_cell mux57 (
    .a (net502),
    .b (net544),
    .sel (net6),
    .out (net545)
  );
  mux_cell mux58 (
    .a (net546),
    .b (net547),
    .sel (net6),
    .out (net548)
  );
  mux_cell mux59 (
    .a (net549),
    .b (net550),
    .sel (net6),
    .out (net551)
  );
  mux_cell mux60 (
    .a (net552),
    .b (net553),
    .sel (net6),
    .out (net554)
  );
  mux_cell mux61 (
    .a (net545),
    .b (net548),
    .sel (net7),
    .out (net555)
  );
  mux_cell mux62 (
    .a (net551),
    .b (net554),
    .sel (net7),
    .out (net556)
  );
  mux_cell mux63 (
    .a (net555),
    .b (net556),
    .sel (net8),
    .out (net36)
  );
  and_cell and143 (
    .a (net529),
    .b (net557),
    .out (net558)
  );
  not_cell not120 (
    .in (net531),
    .out (net557)
  );
  and_cell and144 (
    .a (net559),
    .b (net560),
    .out (net561)
  );
  not_cell not121 (
    .in (net533),
    .out (net559)
  );
  not_cell not122 (
    .in (net535),
    .out (net560)
  );
  and_cell and145 (
    .a (net537),
    .b (net562),
    .out (net563)
  );
  not_cell not123 (
    .in (net539),
    .out (net562)
  );
  not_cell not124 (
    .in (net541),
    .out (net564)
  );
  not_cell not125 (
    .in (net543),
    .out (net565)
  );
  and_cell and146 (
    .a (net564),
    .b (net565),
    .out (net566)
  );
  and_cell and147 (
    .a (net558),
    .b (net561),
    .out (net567)
  );
  and_cell and148 (
    .a (net563),
    .b (net566),
    .out (net568)
  );
  and_cell and149 (
    .a (net567),
    .b (net568),
    .out (net544)
  );
  not_cell not126 (
    .in (net541),
    .out (net569)
  );
  and_cell and150 (
    .a (net570),
    .b (net571),
    .out (net572)
  );
  and_cell and151 (
    .a (net537),
    .b (net539),
    .out (net573)
  );
  and_cell and152 (
    .a (net574),
    .b (net531),
    .out (net575)
  );
  not_cell not127 (
    .in (net533),
    .out (net570)
  );
  not_cell not128 (
    .in (net529),
    .out (net574)
  );
  not_cell not129 (
    .in (net535),
    .out (net571)
  );
  and_cell and153 (
    .a (net569),
    .b (net543),
    .out (net576)
  );
  and_cell and154 (
    .a (net575),
    .b (net572),
    .out (net577)
  );
  and_cell and155 (
    .a (net577),
    .b (net578),
    .out (net546)
  );
  and_cell and156 (
    .a (net573),
    .b (net576),
    .out (net578)
  );
  and_cell and157 (
    .a (net529),
    .b (net531),
    .out (net579)
  );
  and_cell and158 (
    .a (net533),
    .b (net535),
    .out (net580)
  );
  and_cell and159 (
    .a (net537),
    .b (net539),
    .out (net581)
  );
  and_cell and160 (
    .a (net541),
    .b (net582),
    .out (net583)
  );
  and_cell and161 (
    .a (net579),
    .b (net580),
    .out (net584)
  );
  and_cell and162 (
    .a (net581),
    .b (net583),
    .out (net585)
  );
  and_cell and163 (
    .a (net584),
    .b (net585),
    .out (net549)
  );
  not_cell not130 (
    .in (net586),
    .out (net582)
  );
  and_cell and164 (
    .a (net529),
    .b (net535),
    .out (net587)
  );
  and_cell and165 (
    .a (net588),
    .b (net589),
    .out (net590)
  );
  not_cell not131 (
    .in (net531),
    .out (net588)
  );
  not_cell not132 (
    .in (net533),
    .out (net589)
  );
  and_cell and166 (
    .a (net591),
    .b (net592),
    .out (net593)
  );
  not_cell not133 (
    .in (net537),
    .out (net591)
  );
  not_cell not134 (
    .in (net539),
    .out (net592)
  );
  and_cell and167 (
    .a (net541),
    .b (net594),
    .out (net595)
  );
  not_cell not135 (
    .in (net543),
    .out (net594)
  );
  and_cell and168 (
    .a (net595),
    .b (net593),
    .out (net596)
  );
  and_cell and169 (
    .a (net587),
    .b (net590),
    .out (net597)
  );
  and_cell and170 (
    .a (net596),
    .b (net597),
    .out (net550)
  );
  and_cell and171 (
    .a (net529),
    .b (net533),
    .out (net598)
  );
  and_cell and172 (
    .a (net599),
    .b (net600),
    .out (net601)
  );
  and_cell and173 (
    .a (net537),
    .b (net541),
    .out (net602)
  );
  and_cell and174 (
    .a (net603),
    .b (net604),
    .out (net605)
  );
  not_cell not136 (
    .in (net543),
    .out (net604)
  );
  not_cell not137 (
    .in (net539),
    .out (net603)
  );
  not_cell not138 (
    .in (net531),
    .out (net599)
  );
  not_cell not139 (
    .in (net535),
    .out (net600)
  );
  and_cell and175 (
    .a (net598),
    .b (net601),
    .out (net606)
  );
  and_cell and176 (
    .a (net602),
    .b (net605),
    .out (net607)
  );
  and_cell and177 (
    .a (net606),
    .b (net607),
    .out (net552)
  );
  and_cell and178 (
    .a (net530),
    .b (net532),
    .out (net608)
  );
  and_cell and179 (
    .a (net534),
    .b (net536),
    .out (net609)
  );
  and_cell and180 (
    .a (net538),
    .b (net540),
    .out (net610)
  );
  and_cell and181 (
    .a (net542),
    .b (net543),
    .out (net611)
  );
  and_cell and182 (
    .a (net608),
    .b (net609),
    .out (net612)
  );
  and_cell and183 (
    .a (net610),
    .b (net611),
    .out (net613)
  );
  and_cell and184 (
    .a (net612),
    .b (net613),
    .out (net614)
  );
  nand_cell nand1 (
    .a (net612),
    .b (net613),
    .out (net547)
  );
  or_cell or147 (
    .a (net614),
    .b (net547),
    .out (net615)
  );
  or_cell or148 (
    .a (net614),
    .b (net547),
    .out (net616)
  );
  mux_cell mux64 (
    .a (net514),
    .b (net615),
    .sel (net617),
    .out (net52)
  );
  mux_cell mux65 (
    .a (net511),
    .b (net616),
    .sel (net617),
    .out (net68)
  );
  mux_cell mux66 (
    .a (net517),
    .b (net547),
    .sel (net617),
    .out (net84)
  );
  mux_cell mux67 (
    .a (net509),
    .b (net547),
    .sel (net617),
    .out (net100)
  );
  mux_cell mux68 (
    .a (net505),
    .b (net547),
    .sel (net617),
    .out (net116)
  );
  mux_cell mux69 (
    .a (net508),
    .b (net553),
    .sel (net617),
    .out (net132)
  );
endmodule
